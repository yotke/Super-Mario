library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
-- Alex Grinshpun April 2017

entity smileyface_object2 is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer range 0 to 700;
		oCoord_Y	: in integer range 0 to 700;
		ObjectStartX	: in integer range 0 to 700;
		ObjectStartY 	: in integer range 0 to 700;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end smileyface_object2;

architecture behav of smileyface_object2 is 

constant object_X_size : integer := 45;
constant object_Y_size : integer := 56;
constant R_high		: integer := 7;
constant R_low		: integer := 5;
constant G_high		: integer := 4;
constant G_low		: integer := 2;
constant B_high		: integer := 1;
constant B_low		: integer := 0;

type ram_array is array(0 to object_Y_size - 1 , 0 to  object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"F2", x"FF", x"F7", x"F2", x"EE", x"E9", x"E9", x"ED", x"F2", x"F6", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FB", x"F2", x"F2", x"F2", x"F2", x"CD", x"C5", x"C0", x"C5", x"ED", x"F2", x"FB", x"F7", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"FF", x"F2", x"FB", x"F2", x"F2", x"D2", x"FB", x"CD", x"D2", x"F6", x"C0", x"C0", x"C0", x"E9", x"F2", x"F7", x"ED", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"FF", x"FB", x"FB", x"F2", x"CE", x"D6", x"A5", x"A5", x"A9", x"A5", x"FB", x"CD", x"A0", x"C0", x"C0", x"E5", x"EE", x"F6", x"E0", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"FF", x"FF", x"F2", x"A9", x"D6", x"CD", x"CE", x"D2", x"FB", x"A9", x"A9", x"AD", x"A0", x"A0", x"A0", x"C0", x"C5", x"EE", x"F6", x"ED", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"7F", x"F7", x"FB", x"CD", x"80", x"D2", x"C5", x"D6", x"FF", x"FF", x"D6", x"A9", x"84", x"80", x"80", x"A0", x"A0", x"C0", x"C5", x"EE", x"F6", x"F2", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"FF", x"00", x"D2", x"A5", x"80", x"85", x"A9", x"CE", x"D2", x"AD", x"A9", x"85", x"80", x"80", x"80", x"80", x"80", x"A0", x"C0", x"C5", x"EE", x"F7", x"F7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"FB", x"FF", x"AE", x"80", x"80", x"80", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"80", x"80", x"A0", x"C0", x"E9", x"F2", x"E0", x"FB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"D7", x"F7", x"A9", x"60", x"60", x"40", x"40", x"40", x"60", x"60", x"60", x"40", x"40", x"20", x"20", x"40", x"40", x"60", x"80", x"A0", x"C0", x"E9", x"F6", x"F2", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"B2", x"89", x"AE", x"64", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"20", x"20", x"00", x"00", x"00", x"20", x"40", x"60", x"80", x"A0", x"C5", x"EE", x"E5", x"FB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"64", x"89", x"60", x"60", x"40", x"40", x"20", x"00", x"20", x"40", x"40", x"40", x"40", x"20", x"40", x"44", x"20", x"20", x"20", x"20", x"60", x"60", x"A0", x"C9", x"FB", x"F6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"64", x"64", x"60", x"60", x"40", x"20", x"00", x"20", x"20", x"64", x"64", x"88", x"68", x"64", x"68", x"68", x"68", x"64", x"44", x"20", x"20", x"40", x"60", x"A5", x"D2", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"64", x"64", x"60", x"40", x"20", x"20", x"40", x"64", x"64", x"88", x"89", x"89", x"89", x"44", x"49", x"B2", x"8D", x"89", x"89", x"8D", x"44", x"40", x"40", x"80", x"AD", x"A9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"69", x"89", x"60", x"40", x"20", x"44", x"64", x"24", x"8D", x"89", x"A9", x"AD", x"89", x"24", x"05", x"B7", x"D6", x"B1", x"FA", x"FA", x"8D", x"40", x"40", x"60", x"AD", x"89", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"BB", x"89", x"89", x"40", x"40", x"89", x"44", x"05", x"92", x"B2", x"AD", x"AD", x"AD", x"00", x"05", x"BB", x"FF", x"FA", x"FE", x"FF", x"B1", x"64", x"89", x"D6", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"AE", x"B2", x"65", x"65", x"AD", x"44", x"05", x"B7", x"FF", x"FE", x"FE", x"FA", x"6D", x"32", x"DF", x"FF", x"FA", x"FE", x"FE", x"AD", x"64", x"B2", x"F6", x"D1", x"FA", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"DB", x"65", x"89", x"69", x"B1", x"69", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"FF", x"FB", x"DA", x"91", x"DA", x"B6", x"44", x"B1", x"F6", x"FA", x"FA", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"FB", x"FB", x"8E", x"AD", x"B1", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"B2", x"69", x"24", x"6D", x"FF", x"8D", x"B1", x"F6", x"FA", x"FA", x"FA", x"FA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"FF", x"AD", x"D2", x"69", x"8D", x"D2", x"F6", x"FA", x"FE", x"FE", x"FE", x"FE", x"FE", x"D6", x"48", x"24", x"24", x"24", x"69", x"FF", x"DA", x"DA", x"FE", x"FE", x"FE", x"FA", x"FA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"FF", x"84", x"AD", x"69", x"24", x"69", x"B1", x"D2", x"F6", x"F6", x"F6", x"F6", x"F6", x"8D", x"20", x"24", x"20", x"20", x"B1", x"FF", x"FF", x"FF", x"FF", x"FE", x"FA", x"FE", x"FA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"FF", x"AD", x"D2", x"49", x"00", x"00", x"69", x"AD", x"AD", x"B1", x"B1", x"B1", x"8D", x"20", x"20", x"20", x"20", x"8D", x"FA", x"FF", x"FF", x"FA", x"FA", x"FA", x"FA", x"FA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"D6", x"D2", x"F6", x"8D", x"00", x"00", x"00", x"44", x"89", x"89", x"89", x"64", x"20", x"00", x"00", x"20", x"AD", x"FA", x"FA", x"FA", x"FA", x"8D", x"D1", x"D2", x"D1", x"AE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"D6", x"FB", x"5F", x"FB", x"B2", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"64", x"AD", x"FA", x"FA", x"FA", x"F6", x"B1", x"24", x"49", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"FB", x"FB", x"F6", x"D1", x"69", x"44", x"44", x"20", x"24", x"20", x"68", x"AD", x"D1", x"F6", x"F6", x"F6", x"D1", x"AD", x"44", x"20", x"6D", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"FF", x"FF", x"D6", x"D2", x"D1", x"AD", x"AD", x"AD", x"68", x"20", x"D1", x"F6", x"F6", x"F6", x"D1", x"AD", x"89", x"69", x"20", x"20", x"20", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"D6", x"D6", x"B1", x"AD", x"AD", x"8D", x"8D", x"8D", x"B1", x"D6", x"D1", x"D1", x"D1", x"AD", x"64", x"20", x"05", x"2A", x"05", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"FF", x"AD", x"D2", x"64", x"64", x"64", x"64", x"64", x"64", x"89", x"D1", x"D1", x"A9", x"60", x"20", x"20", x"05", x"4F", x"73", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"FF", x"D6", x"FB", x"A9", x"40", x"69", x"8D", x"B6", x"B6", x"B6", x"8D", x"64", x"64", x"40", x"40", x"60", x"60", x"40", x"2A", x"73", x"DB", x"FB", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"FF", x"F7", x"FB", x"AD", x"89", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"44", x"60", x"60", x"80", x"80", x"80", x"80", x"20", x"2E", x"97", x"FF", x"B2", x"D6", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"FB", x"FF", x"AE", x"64", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"4A", x"60", x"80", x"80", x"60", x"60", x"45", x"0A", x"06", x"71", x"FD", x"B5", x"8E", x"92", x"B6", x"FF", x"FF", x"FF", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"FB", x"FF", x"F2", x"A9", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"29", x"25", x"25", x"0A", x"0A", x"0A", x"0F", x"0A", x"29", x"D4", x"D5", x"24", x"8E", x"DB", x"DB", x"DB", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"FF", x"E0", x"F6", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"91", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0F", x"0A", x"25", x"4D", x"24", x"45", x"6E", x"B6", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"FB", x"FB", x"F6", x"F6", x"FF", x"DF", x"DB", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"F8", x"71", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"29", x"00", x"6E", x"DB", x"DB", x"DB", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00"),
(x"FB", x"F2", x"F7", x"EE", x"D2", x"DB", x"DB", x"DB", x"DB", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D5", x"4D", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0F", x"0F", x"0A", x"0A", x"25", x"4E", x"53", x"73", x"77", x"77", x"DB", x"FF", x"FF", x"D6", x"B2", x"AD", x"AD", x"B2", x"DB", x"D7", x"00"),
(x"FB", x"A0", x"D2", x"C9", x"A9", x"DB", x"B7", x"B7", x"B7", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"DB", x"4E", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0B", x"0A", x"0A", x"05", x"06", x"0A", x"0F", x"0F", x"33", x"53", x"73", x"D6", x"B2", x"8D", x"69", x"68", x"69", x"69", x"8D", x"92", x"92"),
(x"FB", x"85", x"AE", x"85", x"84", x"B6", x"96", x"B6", x"B6", x"B7", x"DB", x"DF", x"FF", x"FF", x"DB", x"B6", x"0A", x"0A", x"0B", x"0B", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"06", x"01", x"06", x"06", x"0B", x"0F", x"2F", x"0F", x"4E", x"69", x"64", x"44", x"64", x"8D", x"69", x"44", x"44", x"69", x"FF"),
(x"00", x"AD", x"AE", x"89", x"60", x"8D", x"92", x"96", x"B6", x"92", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"2E", x"0B", x"0B", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"06", x"01", x"06", x"06", x"0B", x"0F", x"0F", x"0A", x"44", x"40", x"40", x"20", x"44", x"8D", x"B1", x"B1", x"8D", x"69", x"69"),
(x"00", x"B6", x"60", x"8D", x"89", x"69", x"92", x"92", x"92", x"92", x"92", x"96", x"DB", x"DB", x"DB", x"72", x"0A", x"0B", x"0B", x"0A", x"0A", x"0A", x"0A", x"0B", x"0B", x"0A", x"06", x"01", x"05", x"06", x"0A", x"0F", x"0A", x"05", x"20", x"20", x"20", x"20", x"89", x"D6", x"F6", x"F5", x"D1", x"AD", x"8D"),
(x"00", x"00", x"FF", x"8D", x"92", x"69", x"92", x"6E", x"6E", x"72", x"6E", x"6D", x"49", x"25", x"05", x"0A", x"0A", x"0F", x"0F", x"0F", x"0B", x"0B", x"0B", x"0B", x"0A", x"0A", x"06", x"01", x"05", x"06", x"0A", x"0B", x"06", x"20", x"20", x"20", x"20", x"44", x"D5", x"F6", x"F6", x"F6", x"D5", x"D1", x"AD"),
(x"00", x"00", x"00", x"00", x"00", x"DF", x"6D", x"72", x"49", x"6E", x"29", x"05", x"01", x"01", x"05", x"0A", x"0F", x"0F", x"0F", x"0F", x"0F", x"0B", x"0A", x"0A", x"0A", x"0A", x"05", x"01", x"05", x"06", x"0A", x"0A", x"01", x"20", x"20", x"20", x"20", x"AD", x"F5", x"FA", x"FA", x"FA", x"F5", x"D1", x"AD"),
(x"00", x"00", x"00", x"00", x"FA", x"FF", x"FF", x"FF", x"BB", x"00", x"2A", x"05", x"05", x"05", x"0A", x"0A", x"0F", x"2F", x"0F", x"0F", x"0B", x"0A", x"0A", x"0A", x"0A", x"06", x"05", x"01", x"05", x"06", x"0A", x"0A", x"01", x"20", x"20", x"00", x"44", x"D1", x"F5", x"FA", x"FA", x"FA", x"F5", x"D1", x"B1"),
(x"00", x"00", x"E8", x"FB", x"FA", x"FF", x"FB", x"B2", x"6D", x"6D", x"4A", x"05", x"05", x"06", x"0A", x"0F", x"2F", x"2F", x"0F", x"0A", x"0A", x"0A", x"06", x"06", x"06", x"06", x"05", x"05", x"05", x"06", x"0A", x"0A", x"00", x"20", x"00", x"00", x"68", x"D1", x"F5", x"FA", x"FA", x"FA", x"F5", x"D1", x"D1"),
(x"00", x"00", x"D6", x"D6", x"D6", x"B6", x"6D", x"45", x"25", x"25", x"4E", x"05", x"06", x"0A", x"0A", x"0F", x"2F", x"0F", x"0A", x"0A", x"06", x"06", x"06", x"05", x"05", x"05", x"05", x"05", x"05", x"06", x"0A", x"0A", x"00", x"20", x"00", x"20", x"8D", x"D1", x"F5", x"FA", x"FA", x"F6", x"D5", x"D1", x"D1"),
(x"00", x"D6", x"F9", x"D6", x"8E", x"49", x"05", x"01", x"01", x"05", x"4A", x"06", x"06", x"0A", x"0B", x"0F", x"0F", x"0A", x"0A", x"06", x"06", x"05", x"05", x"05", x"05", x"05", x"09", x"29", x"2A", x"0A", x"0A", x"05", x"20", x"20", x"00", x"20", x"8D", x"D1", x"D1", x"D5", x"D5", x"D5", x"D1", x"D1", x"B1"),
(x"00", x"D6", x"D6", x"92", x"49", x"05", x"05", x"06", x"2A", x"4E", x"2A", x"06", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"06", x"05", x"05", x"05", x"29", x"29", x"4A", x"4A", x"4E", x"6E", x"2A", x"0A", x"05", x"20", x"20", x"00", x"40", x"88", x"8D", x"8D", x"AD", x"AD", x"B1", x"B1", x"B1", x"B1"),
(x"FB", x"00", x"B2", x"49", x"06", x"06", x"0A", x"2A", x"2A", x"4E", x"0A", x"06", x"0A", x"0A", x"0A", x"0A", x"0A", x"06", x"06", x"06", x"06", x"05", x"29", x"4E", x"92", x"6E", x"00", x"B6", x"4E", x"6E", x"2A", x"00", x"20", x"20", x"20", x"64", x"68", x"68", x"68", x"88", x"89", x"8D", x"AD", x"88", x"AD"),
(x"B2", x"B6", x"6D", x"25", x"0A", x"0A", x"0A", x"0A", x"2E", x"2E", x"06", x"0A", x"0A", x"0A", x"0A", x"06", x"06", x"06", x"06", x"06", x"0A", x"2A", x"6E", x"4E", x"00", x"00", x"00", x"00", x"6E", x"73", x"05", x"20", x"20", x"20", x"20", x"8D", x"AD", x"AD", x"B1", x"AD", x"AD", x"AD", x"D1", x"B1", x"00"),
(x"D2", x"8E", x"44", x"05", x"0A", x"0A", x"0A", x"0A", x"4E", x"0A", x"06", x"0A", x"0A", x"0A", x"06", x"06", x"06", x"06", x"06", x"0A", x"2A", x"4E", x"4E", x"DB", x"00", x"00", x"00", x"00", x"2A", x"53", x"05", x"24", x"20", x"20", x"68", x"AD", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"00"),
(x"B2", x"69", x"20", x"05", x"0A", x"0A", x"2E", x"2E", x"4F", x"0A", x"06", x"06", x"0A", x"0A", x"06", x"06", x"06", x"06", x"0A", x"2A", x"6E", x"2A", x"B6", x"00", x"00", x"00", x"00", x"00", x"4E", x"00", x"29", x"24", x"20", x"20", x"88", x"D1", x"D1", x"F5", x"D5", x"D1", x"D1", x"B1", x"B1", x"00", x"00"),
(x"6D", x"44", x"20", x"05", x"06", x"0A", x"2E", x"4F", x"2F", x"0A", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"0A", x"2A", x"6E", x"06", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2A", x"2A", x"49", x"24", x"44", x"AD", x"D1", x"D5", x"F6", x"D5", x"D1", x"B1", x"B1", x"B1", x"00", x"00"),
(x"49", x"20", x"00", x"01", x"05", x"0A", x"2A", x"2F", x"2E", x"0A", x"0A", x"06", x"06", x"06", x"06", x"0A", x"0A", x"2A", x"4E", x"00", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"6D", x"6D", x"44", x"44", x"AD", x"D1", x"D1", x"D1", x"D1", x"AD", x"88", x"AD", x"00", x"00", x"00"),
(x"44", x"20", x"20", x"00", x"05", x"06", x"2A", x"2E", x"2A", x"0A", x"0A", x"0A", x"0A", x"06", x"0A", x"0A", x"2A", x"4E", x"FF", x"72", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"6D", x"49", x"8D", x"B1", x"D1", x"B1", x"AD", x"88", x"AD", x"00", x"00", x"00", x"00"),
(x"20", x"20", x"20", x"20", x"00", x"05", x"4E", x"4E", x"2A", x"2A", x"0A", x"0A", x"0A", x"0A", x"0A", x"2A", x"4E", x"FF", x"72", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"68", x"44", x"AD", x"AD", x"88", x"AD", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"20", x"20", x"20", x"20", x"20", x"24", x"49", x"6E", x"4E", x"2A", x"2A", x"2A", x"0A", x"2A", x"2A", x"4E", x"01", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"44", x"20", x"20", x"20", x"20", x"20", x"44", x"69", x"92", x"6E", x"4E", x"4E", x"4A", x"4E", x"6E", x"4E", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"20", x"24", x"20", x"20", x"44", x"44", x"68", x"6D", x"69", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("000000111111111111100000000000000000000000000"),
("000001111111111111111000000000000000000000000"),
("000011111111111111111100000000000000000000000"),
("000111111111111111111110000000000000000000000"),
("000111111111111111111111000000000000000000000"),
("001111111111111111111111100000000000000000000"),
("001011111111111111111111100000000000000000000"),
("001111111111111111111111110000000000000000000"),
("001111111111111111111111110000000000000000000"),
("011111111111111000111111111000000000000000000"),
("011111110111111111111111111000000000000000000"),
("011111101111111111111111111000000000000000000"),
("011111111111111111111111111000000000000000000"),
("011111111111111111111111111100000000000000000"),
("011111111111110111111111111110000000000000000"),
("001111111111111111111111111110000000000000000"),
("001111111111111111111111111110000000000000000"),
("000111111111111111111111111110000000000000000"),
("001111111111111111111111111110000000000000000"),
("001111111111111111111111111110000000000000000"),
("001111001111111111111111111100000000000000000"),
("001111000111111001111111111100000000000000000"),
("001111110000000111111111110000000000000000000"),
("000011111111111111111111110000000000000000000"),
("000011111111111111111111110000000000000000000"),
("000001111111111111111111111111110000000000000"),
("000001111111111111111111111111111000000000000"),
("000011111111111111111111111111111100000000000"),
("000111111111111111111111111111111100000000000"),
("000111111111111111111111111111111110000000000"),
("001111111111111111111111111111111110000000000"),
("011111111111111111111111111111111110000000000"),
("011111111111111111111111111101111110111111000"),
("111111111111111111111111111111111111111111110"),
("111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111"),
("000001111111111111111111111111111111111111111"),
("000011111011111111111111111111111110111111111"),
("001111111111111111111111111111110100111111111"),
("001111111111111111111111111111110101111111111"),
("011111111111111111111111111111111101111111111"),
("011111111111111111111111111111111101111111111"),
("101111111111111111111111110111101111111111111"),
("111111111111111111111111000011111111111111110"),
("111111111111111111111111000011111111111111110"),
("111111111111111111111110000010111111111111100"),
("111111111111111111111100000001111111111111100"),
("110111111111111111101000000001111111111111000"),
("111011111111111111110000000000011111111110000"),
("111101111111111111100000000000000111111000000"),
("111111111111111111000000000000000000000000000"),
("111111111111111110000000000000000000000000000"),
("111111111111110000000000000000000000000000000")
);



signal bCoord_X : integer := 0;
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--		
signal objectWestXboundary : integer;
signal objectSouthboundary : integer;
signal objectXboundariesTrue : boolean;
signal objectYboundariesTrue : boolean;
signal ObjectStartX_d : integer;
--signal keepflag : std_logic;
attribute syn_keep: boolean;
--attribute syn_keep of keepflag: signal is true;
attribute preserve : boolean;
--attribute preserve of keepflag: signal is true;
attribute noprune: boolean;  
--attribute noprune of keepflag: signal is true;
begin

-- Calculate object boundaries
objectWestXboundary	<= object_X_size+ObjectStartX;
objectSouthboundary	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectWestXboundary) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectSouthboundary) else '0';

	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)

  		
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;
		ObjectStartX_d <= 0;

		elsif CLK'event and CLK='1' then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
			ObjectStartX_d <= ObjectStartX;
	end if;

  end process;

	--keepflag <= '1' when 	ObjectStartX - ObjectStartX_d > 100 else '0';	
		
end behav;		
		