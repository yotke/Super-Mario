--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bombTableTC is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(12 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end bombTableTC;

architecture arch of bombTableTC is

type table_type is array(0 to 8191) of std_logic_vector(7 downto 0);
signal sin_table : table_type;

begin

  SinTableTC_proc: process(RESET_N, CLK)
    constant sin_table : table_type := (
X"00",
X"06",
X"0C",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"07",
X"06",
X"06",
X"06",
X"06",
X"05",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"01",
X"FB",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"00",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"FA",
X"F5",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"F9",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"01",
X"03",
X"FE",
X"F5",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"05",
X"09",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FA",
X"F6",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FA",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"04",
X"0A",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"FE",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FF",
X"06",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"F9",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"05",
X"0A",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"F6",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"04",
X"0A",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FA",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FD",
X"01",
X"0A",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"FE",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"02",
X"0A",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"F7",
X"F5",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"04",
X"0A",
X"08",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"FC",
X"F5",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"02",
X"0A",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"F7",
X"F5",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FD",
X"00",
X"0A",
X"08",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"03",
X"0A",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"FF",
X"F5",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"01",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"01",
X"06",
X"04",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"F7",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FA",
X"FD",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"00",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"04",
X"07",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"04",
X"00",
X"F7",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FE",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"05",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"04",
X"03",
X"04",
X"00",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"04",
X"08",
X"06",
X"07",
X"05",
X"06",
X"05",
X"06",
X"05",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"F9",
X"F7",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"02",
X"08",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"FC",
X"F8",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"00",
X"08",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FC",
X"F7",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"FE",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"FB",
X"F7",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"00",
X"08",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"03",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"04",
X"03",
X"04",
X"02",
X"04",
X"00",
X"F7",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"05",
X"08",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"FB",
X"F7",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"04",
X"08",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"02",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"00",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FA",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"07",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FD",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"09",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FB",
X"F6",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"04",
X"08",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"01",
X"FA",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"04",
X"08",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"03",
X"01",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"00",
X"06",
X"08",
X"07",
X"07",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"03",
X"FC",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"05",
X"09",
X"07",
X"08",
X"07",
X"07",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FA",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"00",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"FC",
X"F6",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FF",
X"05",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"FE",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FF",
X"08",
X"08",
X"07",
X"08",
X"07",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"04",
X"09",
X"08",
X"08",
X"07",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FB",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"01",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"01",
X"02",
X"01",
X"02",
X"FF",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"05",
X"0A",
X"08",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"F8",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"02",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"F8",
X"F5",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"02",
X"FF",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"03",
X"0A",
X"08",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"F7",
X"F5",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"02",
X"0B",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"F9",
X"F4",
X"F7",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"09",
X"0B",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"F8",
X"F4",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"04",
X"0B",
X"09",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"F9",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FA",
X"F3",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"09",
X"0C",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"07",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00"






  );
  begin

    if (RESET_N='0') then
      Q <= sin_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sin_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;