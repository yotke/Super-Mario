--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity obstacleTableTC is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(12 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end obstacleTableTC;

architecture arch of obstacleTableTC is

type table_type is array(0 to 8191) of std_logic_vector(7 downto 0);
signal sin_table : table_type;

begin

  SinTableTC_proc: process(RESET_N, CLK)
    constant sin_table : table_type := (
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"02",
X"08",
X"08",
X"04",
X"FB",
X"F2",
X"F2",
X"F4",
X"F5",
X"F8",
X"FA",
X"F7",
X"F8",
X"FB",
X"FA",
X"FA",
X"FC",
X"FD",
X"00",
X"0B",
X"15",
X"10",
X"0D",
X"0E",
X"11",
X"0E",
X"09",
X"0D",
X"06",
X"00",
X"00",
X"04",
X"01",
X"F7",
X"F7",
X"F6",
X"F7",
X"F1",
X"EE",
X"F0",
X"F1",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F5",
X"F7",
X"F8",
X"FD",
X"05",
X"0D",
X"13",
X"15",
X"12",
X"0F",
X"0F",
X"0E",
X"0D",
X"0F",
X"10",
X"0F",
X"10",
X"10",
X"0E",
X"0D",
X"0D",
X"0D",
X"05",
X"FA",
X"F1",
X"EE",
X"EE",
X"EE",
X"F0",
X"F0",
X"F0",
X"F1",
X"F0",
X"F0",
X"F1",
X"F3",
X"F5",
X"F5",
X"F8",
X"FC",
X"00",
X"0A",
X"0F",
X"0F",
X"12",
X"12",
X"10",
X"10",
X"11",
X"0F",
X"0D",
X"0D",
X"0D",
X"0B",
X"07",
X"00",
X"F9",
X"F5",
X"FB",
X"F8",
X"F1",
X"F6",
X"F7",
X"F1",
X"EE",
X"F0",
X"F1",
X"F1",
X"F1",
X"F4",
X"F6",
X"F9",
X"F7",
X"FA",
X"00",
X"00",
X"0C",
X"12",
X"0E",
X"11",
X"12",
X"12",
X"10",
X"0F",
X"10",
X"10",
X"0F",
X"0F",
X"0E",
X"0D",
X"0C",
X"0C",
X"0C",
X"09",
X"08",
X"03",
X"F8",
X"EF",
X"EB",
X"EB",
X"EB",
X"EC",
X"ED",
X"F2",
X"F4",
X"F1",
X"EF",
X"F1",
X"F2",
X"F1",
X"F1",
X"F1",
X"F0",
X"F2",
X"FD",
X"04",
X"09",
X"0E",
X"0F",
X"12",
X"13",
X"12",
X"11",
X"11",
X"10",
X"0F",
X"0E",
X"0E",
X"0F",
X"0D",
X"0C",
X"08",
X"05",
X"00",
X"FA",
X"F4",
X"EE",
X"EC",
X"ED",
X"EE",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"F0",
X"F2",
X"F5",
X"FA",
X"FB",
X"00",
X"03",
X"08",
X"0E",
X"0F",
X"11",
X"10",
X"10",
X"10",
X"0D",
X"0D",
X"0F",
X"0D",
X"0B",
X"0C",
X"0A",
X"05",
X"02",
X"01",
X"00",
X"F9",
X"F0",
X"EB",
X"EB",
X"ED",
X"EE",
X"EE",
X"ED",
X"ED",
X"EE",
X"EE",
X"EF",
X"F0",
X"F0",
X"F3",
X"F5",
X"F6",
X"F9",
X"FA",
X"FF",
X"04",
X"04",
X"04",
X"0A",
X"0B",
X"0F",
X"12",
X"11",
X"11",
X"11",
X"0F",
X"0E",
X"0E",
X"0D",
X"0B",
X"0A",
X"07",
X"07",
X"09",
X"07",
X"04",
X"02",
X"00",
X"FC",
X"FE",
X"01",
X"00",
X"00",
X"02",
X"01",
X"FF",
X"FE",
X"FD",
X"FC",
X"FA",
X"FA",
X"FC",
X"FD",
X"F9",
X"F8",
X"FE",
X"FA",
X"F5",
X"F2",
X"F2",
X"F8",
X"F8",
X"FB",
X"FC",
X"F7",
X"F3",
X"F0",
X"F0",
X"F3",
X"F5",
X"F5",
X"FA",
X"FB",
X"FA",
X"F9",
X"F8",
X"F7",
X"F7",
X"F8",
X"FC",
X"00",
X"01",
X"04",
X"06",
X"08",
X"01",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"04",
X"07",
X"09",
X"07",
X"07",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0B",
X"0A",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0B",
X"0A",
X"06",
X"05",
X"04",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FD",
X"FC",
X"FA",
X"FA",
X"FC",
X"FA",
X"F4",
X"F1",
X"F3",
X"F5",
X"F4",
X"F2",
X"F3",
X"F6",
X"F7",
X"F9",
X"F9",
X"F6",
X"F3",
X"F3",
X"F4",
X"F7",
X"F7",
X"F7",
X"FA",
X"FB",
X"FE",
X"00",
X"00",
X"02",
X"06",
X"05",
X"04",
X"06",
X"06",
X"02",
X"FF",
X"FB",
X"FA",
X"FD",
X"00",
X"03",
X"04",
X"06",
X"08",
X"0D",
X"0F",
X"0E",
X"0D",
X"0C",
X"09",
X"04",
X"04",
X"06",
X"05",
X"02",
X"00",
X"00",
X"FE",
X"FA",
X"FC",
X"03",
X"0B",
X"0C",
X"0B",
X"09",
X"08",
X"05",
X"04",
X"04",
X"02",
X"03",
X"01",
X"00",
X"00",
X"01",
X"03",
X"03",
X"01",
X"FD",
X"FB",
X"FC",
X"FB",
X"F7",
X"F6",
X"FA",
X"00",
X"00",
X"01",
X"02",
X"00",
X"FD",
X"F9",
X"F6",
X"F6",
X"F6",
X"F5",
X"F6",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FB",
X"F8",
X"F7",
X"F8",
X"FB",
X"FE",
X"FF",
X"04",
X"0E",
X"11",
X"0E",
X"0C",
X"0D",
X"0D",
X"0B",
X"0B",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0A",
X"07",
X"04",
X"01",
X"00",
X"FD",
X"FA",
X"F9",
X"FB",
X"FB",
X"F7",
X"F5",
X"F6",
X"F6",
X"F7",
X"FC",
X"FA",
X"F8",
X"FE",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"00",
X"00",
X"00",
X"00",
X"04",
X"0C",
X"0E",
X"0E",
X"0D",
X"0C",
X"0C",
X"0B",
X"0B",
X"07",
X"00",
X"FC",
X"F9",
X"F8",
X"F7",
X"F4",
X"F2",
X"F1",
X"F4",
X"F5",
X"F5",
X"F4",
X"F3",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F5",
X"F5",
X"F5",
X"F7",
X"F8",
X"F9",
X"FA",
X"FC",
X"FC",
X"FB",
X"F9",
X"FA",
X"FC",
X"FF",
X"00",
X"00",
X"00",
X"03",
X"07",
X"0A",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"09",
X"09",
X"08",
X"07",
X"07",
X"06",
X"04",
X"01",
X"FF",
X"FE",
X"00",
X"02",
X"03",
X"04",
X"07",
X"07",
X"06",
X"06",
X"08",
X"09",
X"08",
X"06",
X"05",
X"02",
X"00",
X"00",
X"00",
X"01",
X"02",
X"00",
X"FF",
X"00",
X"02",
X"02",
X"00",
X"FC",
X"FB",
X"FC",
X"FC",
X"FB",
X"FB",
X"FA",
X"FA",
X"FB",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"F9",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F5",
X"F3",
X"F4",
X"F4",
X"F3",
X"F4",
X"F6",
X"F7",
X"FA",
X"FC",
X"FE",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"02",
X"05",
X"08",
X"09",
X"09",
X"07",
X"08",
X"0B",
X"0D",
X"0A",
X"0A",
X"0A",
X"09",
X"06",
X"01",
X"01",
X"02",
X"00",
X"00",
X"01",
X"02",
X"04",
X"05",
X"05",
X"07",
X"08",
X"08",
X"07",
X"05",
X"06",
X"07",
X"05",
X"03",
X"00",
X"00",
X"01",
X"02",
X"02",
X"03",
X"04",
X"06",
X"07",
X"08",
X"07",
X"05",
X"05",
X"04",
X"03",
X"01",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FE",
X"FB",
X"F6",
X"F5",
X"F6",
X"F6",
X"F3",
X"F0",
X"EE",
X"EC",
X"EC",
X"EB",
X"ED",
X"ED",
X"EE",
X"F0",
X"F2",
X"F2",
X"F1",
X"F1",
X"F2",
X"F3",
X"F4",
X"F6",
X"F9",
X"FC",
X"FD",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"04",
X"07",
X"09",
X"08",
X"07",
X"08",
X"0A",
X"0A",
X"09",
X"07",
X"06",
X"07",
X"07",
X"04",
X"02",
X"00",
X"00",
X"01",
X"04",
X"07",
X"08",
X"08",
X"07",
X"08",
X"09",
X"09",
X"08",
X"08",
X"08",
X"06",
X"05",
X"04",
X"03",
X"01",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"02",
X"03",
X"03",
X"01",
X"02",
X"03",
X"06",
X"04",
X"02",
X"00",
X"00",
X"00",
X"FF",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FA",
X"FA",
X"F7",
X"F2",
X"F2",
X"F3",
X"F4",
X"F4",
X"F3",
X"F4",
X"F4",
X"F3",
X"F4",
X"F5",
X"F5",
X"F5",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F9",
X"FC",
X"FD",
X"FE",
X"FC",
X"FC",
X"FD",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"03",
X"05",
X"08",
X"0A",
X"09",
X"0A",
X"09",
X"07",
X"06",
X"05",
X"07",
X"09",
X"0B",
X"09",
X"07",
X"07",
X"08",
X"08",
X"07",
X"05",
X"04",
X"03",
X"02",
X"01",
X"00",
X"00",
X"FE",
X"FD",
X"FE",
X"FF",
X"FF",
X"FE",
X"FD",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"05",
X"07",
X"07",
X"06",
X"05",
X"05",
X"05",
X"06",
X"06",
X"04",
X"03",
X"02",
X"02",
X"02",
X"01",
X"00",
X"01",
X"02",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FD",
X"FC",
X"FC",
X"FD",
X"00",
X"00",
X"FE",
X"FA",
X"F8",
X"F9",
X"FA",
X"FD",
X"00",
X"FD",
X"F9",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F7",
X"F7",
X"F8",
X"F8",
X"F7",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F8",
X"FA",
X"FA",
X"F9",
X"FA",
X"FB",
X"FA",
X"FB",
X"FD",
X"FE",
X"FE",
X"FD",
X"FC",
X"FD",
X"FF",
X"FF",
X"FE",
X"FE",
X"FF",
X"00",
X"01",
X"03",
X"06",
X"08",
X"09",
X"09",
X"08",
X"08",
X"0A",
X"0B",
X"0C",
X"0B",
X"0A",
X"0A",
X"0C",
X"0D",
X"0F",
X"0F",
X"0F",
X"0E",
X"0D",
X"0C",
X"0C",
X"0B",
X"0B",
X"0A",
X"0A",
X"09",
X"07",
X"06",
X"05",
X"04",
X"05",
X"05",
X"04",
X"03",
X"04",
X"04",
X"03",
X"02",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"FD",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"F9",
X"F7",
X"F6",
X"F5",
X"F5",
X"F4",
X"F3",
X"F2",
X"F2",
X"F2",
X"F2",
X"F1",
X"F2",
X"F2",
X"F3",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F4",
X"F6",
X"F8",
X"F8",
X"F7",
X"F7",
X"F7",
X"F9",
X"FA",
X"FB",
X"FC",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"02",
X"03",
X"03",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"03",
X"04",
X"04",
X"03",
X"03",
X"04",
X"05",
X"07",
X"09",
X"0C",
X"0D",
X"0D",
X"0D",
X"0D",
X"0E",
X"0F",
X"0F",
X"0E",
X"0D",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"09",
X"08",
X"07",
X"04",
X"01",
X"00",
X"FF",
X"FE",
X"FC",
X"FB",
X"FA",
X"FB",
X"FC",
X"FD",
X"FE",
X"FE",
X"FE",
X"FC",
X"FA",
X"F9",
X"FA",
X"FB",
X"FD",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"04",
X"05",
X"06",
X"07",
X"08",
X"07",
X"05",
X"03",
X"03",
X"03",
X"04",
X"03",
X"02",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FD",
X"FA",
X"F8",
X"F8",
X"FA",
X"FB",
X"FB",
X"FA",
X"F8",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F5",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F8",
X"FA",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"00",
X"00",
X"01",
X"02",
X"04",
X"05",
X"06",
X"07",
X"08",
X"0B",
X"0C",
X"0E",
X"0F",
X"0F",
X"0F",
X"0E",
X"0D",
X"0B",
X"0B",
X"0B",
X"0A",
X"09",
X"08",
X"08",
X"08",
X"07",
X"07",
X"08",
X"08",
X"08",
X"07",
X"06",
X"06",
X"04",
X"03",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"02",
X"03",
X"03",
X"02",
X"03",
X"03",
X"04",
X"05",
X"06",
X"05",
X"04",
X"03",
X"03",
X"02",
X"01",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"F9",
X"F9",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F6",
X"F6",
X"F4",
X"F2",
X"F1",
X"F1",
X"F1",
X"F0",
X"F0",
X"F0",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F2",
X"F4",
X"F5",
X"F6",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"03",
X"04",
X"06",
X"06",
X"05",
X"04",
X"03",
X"04",
X"05",
X"07",
X"09",
X"0A",
X"09",
X"07",
X"08",
X"09",
X"0A",
X"0C",
X"0C",
X"0C",
X"0B",
X"0A",
X"08",
X"08",
X"07",
X"07",
X"07",
X"06",
X"06",
X"05",
X"04",
X"03",
X"02",
X"02",
X"03",
X"04",
X"04",
X"04",
X"03",
X"03",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FB",
X"F9",
X"F7",
X"F7",
X"F7",
X"F8",
X"F9",
X"FA",
X"FC",
X"FE",
X"00",
X"01",
X"02",
X"03",
X"03",
X"04",
X"04",
X"05",
X"05",
X"05",
X"04",
X"06",
X"07",
X"08",
X"07",
X"06",
X"06",
X"06",
X"07",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"06",
X"06",
X"07",
X"07",
X"07",
X"06",
X"05",
X"03",
X"03",
X"02",
X"01",
X"01",
X"00",
X"00",
X"FE",
X"FB",
X"FA",
X"F9",
X"F7",
X"F7",
X"F6",
X"F5",
X"F4",
X"F4",
X"F3",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F2",
X"F3",
X"F3",
X"F3",
X"F4",
X"F5",
X"F4",
X"F3",
X"F3",
X"F3",
X"F2",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F3",
X"F2",
X"F2",
X"F1",
X"F1",
X"F2",
X"F3",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F7",
X"F8",
X"F9",
X"FB",
X"FD",
X"FF",
X"00",
X"00",
X"02",
X"03",
X"05",
X"05",
X"06",
X"08",
X"09",
X"09",
X"0A",
X"0B",
X"0C",
X"0B",
X"0B",
X"0B",
X"0C",
X"0C",
X"0C",
X"0D",
X"0C",
X"0C",
X"0B",
X"0A",
X"09",
X"08",
X"07",
X"07",
X"07",
X"08",
X"09",
X"09",
X"09",
X"08",
X"07",
X"06",
X"06",
X"05",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"03",
X"03",
X"05",
X"06",
X"08",
X"08",
X"08",
X"07",
X"05",
X"05",
X"04",
X"04",
X"04",
X"03",
X"03",
X"02",
X"02",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FE",
X"FE",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FD",
X"FB",
X"FB",
X"FB",
X"FB",
X"FA",
X"F9",
X"F8",
X"F7",
X"F6",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F7",
X"F7",
X"F6",
X"F5",
X"F5",
X"F5",
X"F6",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FB",
X"FD",
X"FE",
X"00",
X"00",
X"00",
X"01",
X"02",
X"03",
X"03",
X"02",
X"02",
X"02",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"02",
X"02",
X"04",
X"06",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"08",
X"09",
X"09",
X"09",
X"08",
X"07",
X"06",
X"06",
X"06",
X"06",
X"07",
X"07",
X"07",
X"08",
X"09",
X"09",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"08",
X"08",
X"07",
X"06",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FC",
X"FB",
X"FA",
X"FA",
X"FA",
X"FB",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FD",
X"FC",
X"FC",
X"FB",
X"FB",
X"F9",
X"F8",
X"F7",
X"F7",
X"F7",
X"F7",
X"F6",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F4",
X"F4",
X"F5",
X"F6",
X"F7",
X"F8",
X"F9",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FE",
X"FE",
X"FF",
X"FE",
X"FD",
X"FC",
X"FB",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FC",
X"FC",
X"FB",
X"FB",
X"FA",
X"FA",
X"F9",
X"F9",
X"F8",
X"F9",
X"F9",
X"FB",
X"FC",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"02",
X"02",
X"03",
X"05",
X"05",
X"05",
X"05",
X"06",
X"05",
X"06",
X"07",
X"08",
X"09",
X"0A",
X"0B",
X"0C",
X"0D",
X"0D",
X"0E",
X"0E",
X"0E",
X"0E",
X"0E",
X"0E",
X"0E",
X"0F",
X"10",
X"11",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0D",
X"0C",
X"0B",
X"0B",
X"0A",
X"09",
X"08",
X"06",
X"05",
X"04",
X"03",
X"03",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FC",
X"FB",
X"F9",
X"F8",
X"F8",
X"F7",
X"F6",
X"F6",
X"F5",
X"F4",
X"F4",
X"F4",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F5",
X"F6",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"FA",
X"FB",
X"FC",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"FB",
X"FB",
X"FA",
X"FA",
X"F9",
X"F9",
X"F9",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"FA",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"02",
X"04",
X"06",
X"07",
X"08",
X"08",
X"08",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"07",
X"08",
X"09",
X"0A",
X"0C",
X"0C",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"08",
X"07",
X"06",
X"05",
X"05",
X"04",
X"03",
X"03",
X"02",
X"02",
X"02",
X"03",
X"03",
X"04",
X"04",
X"04",
X"04",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"03",
X"02",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FB",
X"FA",
X"FA",
X"FA",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FC",
X"FD",
X"FE",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FC",
X"FB",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"F9",
X"F8",
X"F7",
X"F6",
X"F6",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F8",
X"F9",
X"FB",
X"FC",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"02",
X"04",
X"05",
X"06",
X"08",
X"08",
X"09",
X"0A",
X"0A",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"05",
X"04",
X"03",
X"02",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"FE",
X"FD",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"02",
X"04",
X"05",
X"07",
X"07",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"06",
X"06",
X"05",
X"04",
X"04",
X"03",
X"03",
X"03",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"FE",
X"FC",
X"FA",
X"F9",
X"F8",
X"F7",
X"F6",
X"F5",
X"F4",
X"F2",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F1",
X"F1",
X"F0",
X"F0",
X"F0",
X"EF",
X"EF",
X"EF",
X"F0",
X"F1",
X"F2",
X"F3",
X"F4",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F5",
X"F6",
X"F7",
X"F9",
X"FA",
X"FD",
X"FF",
X"00",
X"01",
X"02",
X"03",
X"03",
X"05",
X"06",
X"07",
X"07",
X"07",
X"07",
X"07",
X"08",
X"08",
X"08",
X"08",
X"08",
X"09",
X"09",
X"09",
X"07",
X"06",
X"05",
X"04",
X"05",
X"05",
X"05",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"05",
X"04",
X"03",
X"04",
X"06",
X"07",
X"08",
X"08",
X"07",
X"07",
X"07",
X"08",
X"08",
X"08",
X"07",
X"07",
X"06",
X"06",
X"05",
X"04",
X"03",
X"02",
X"02",
X"02",
X"02",
X"03",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FC",
X"FA",
X"F9",
X"F8",
X"F7",
X"F6",
X"F5",
X"F4",
X"F3",
X"F2",
X"F2",
X"F2",
X"F2",
X"F1",
X"F1",
X"F1",
X"F1",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F3",
X"F4",
X"F5",
X"F5",
X"F4",
X"F5",
X"F7",
X"F8",
X"F9",
X"F9",
X"FA",
X"FA",
X"FC",
X"FE",
X"00",
X"00",
X"01",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"02",
X"04",
X"06",
X"07",
X"07",
X"07",
X"07",
X"08",
X"09",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"0B",
X"0C",
X"0D",
X"0D",
X"0D",
X"0C",
X"0B",
X"09",
X"07",
X"07",
X"07",
X"07",
X"06",
X"05",
X"03",
X"01",
X"02",
X"02",
X"00",
X"FF",
X"FE",
X"FF",
X"FF",
X"FC",
X"F8",
X"F5",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F6",
X"F7",
X"FA",
X"FC",
X"FD",
X"FD",
X"FF",
X"00",
X"02",
X"02",
X"01",
X"01",
X"00",
X"FF",
X"FD",
X"FE",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"02",
X"02",
X"03",
X"03",
X"02",
X"01",
X"02",
X"02",
X"02",
X"02",
X"04",
X"06",
X"08",
X"08",
X"09",
X"0A",
X"0A",
X"0A",
X"09",
X"08",
X"07",
X"05",
X"03",
X"02",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FD",
X"FB",
X"FA",
X"F9",
X"F9",
X"FA",
X"FB",
X"FA",
X"FA",
X"F8",
X"F5",
X"F0",
X"ED",
X"EE",
X"EE",
X"EF",
X"EF",
X"F0",
X"F1",
X"F2",
X"F3",
X"F3",
X"F5",
X"F5",
X"F5",
X"F6",
X"F9",
X"FB",
X"FD",
X"FE",
X"FF",
X"00",
X"02",
X"04",
X"06",
X"07",
X"09",
X"0C",
X"0D",
X"0E",
X"0D",
X"0C",
X"0B",
X"0B",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"0C",
X"0A",
X"07",
X"06",
X"04",
X"02",
X"00",
X"00",
X"01",
X"02",
X"02",
X"01",
X"00",
X"00",
X"01",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"02",
X"03",
X"03",
X"04",
X"04",
X"03",
X"02",
X"00",
X"FD",
X"FB",
X"FB",
X"FA",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FB",
X"FC",
X"FD",
X"FD",
X"FE",
X"00",
X"00",
X"02",
X"04",
X"05",
X"07",
X"09",
X"0B",
X"0A",
X"07",
X"05",
X"03",
X"01",
X"01",
X"02",
X"02",
X"03",
X"04",
X"03",
X"01",
X"00",
X"FF",
X"FE",
X"FC",
X"FC",
X"FB",
X"FC",
X"FB",
X"F9",
X"F6",
X"F4",
X"F3",
X"F1",
X"EE",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EF",
X"F1",
X"F5",
X"FA",
X"FD",
X"FF",
X"00",
X"00",
X"01",
X"04",
X"06",
X"06",
X"06",
X"06",
X"04",
X"04",
X"01",
X"00",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"02",
X"05",
X"06",
X"08",
X"09",
X"08",
X"07",
X"07",
X"04",
X"00",
X"FF",
X"FF",
X"FD",
X"FA",
X"F8",
X"F7",
X"F7",
X"F6",
X"F6",
X"F7",
X"F9",
X"FA",
X"FC",
X"FE",
X"00",
X"00",
X"00",
X"01",
X"03",
X"05",
X"05",
X"06",
X"06",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"02",
X"02",
X"02",
X"03",
X"05",
X"06",
X"08",
X"08",
X"08",
X"07",
X"05",
X"02",
X"00",
X"00",
X"FF",
X"FE",
X"FC",
X"FB",
X"F9",
X"F9",
X"FA",
X"FA",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"FB",
X"FC",
X"FD",
X"FD",
X"FF",
X"01",
X"03",
X"05",
X"05",
X"04",
X"04",
X"05",
X"05",
X"05",
X"04",
X"02",
X"00",
X"00",
X"04",
X"08",
X"08",
X"06",
X"02",
X"FF",
X"FE",
X"FD",
X"FE",
X"FE",
X"FA",
X"F6",
X"F6",
X"F5",
X"F2",
X"F1",
X"F3",
X"F5",
X"F8",
X"F9",
X"FA",
X"F9",
X"F9",
X"FB",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"03",
X"05",
X"05",
X"04",
X"04",
X"03",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"F9",
X"F8",
X"F7",
X"F4",
X"F3",
X"F3",
X"F4",
X"F6",
X"F8",
X"F9",
X"F9",
X"FD",
X"00",
X"03",
X"07",
X"0B",
X"0D",
X"0B",
X"09",
X"07",
X"04",
X"02",
X"01",
X"02",
X"04",
X"06",
X"04",
X"01",
X"00",
X"01",
X"03",
X"04",
X"01",
X"FE",
X"FC",
X"F9",
X"F7",
X"F5",
X"F4",
X"F6",
X"FA",
X"FD",
X"00",
X"02",
X"04",
X"04",
X"05",
X"07",
X"08",
X"07",
X"06",
X"09",
X"0B",
X"0C",
X"0C",
X"0B",
X"0A",
X"09",
X"08",
X"06",
X"03",
X"00",
X"FD",
X"F9",
X"F7",
X"F7",
X"F7",
X"F8",
X"FB",
X"FD",
X"00",
X"03",
X"03",
X"05",
X"09",
X"0A",
X"0A",
X"06",
X"03",
X"04",
X"03",
X"01",
X"00",
X"00",
X"02",
X"05",
X"06",
X"06",
X"07",
X"05",
X"01",
X"FC",
X"FC",
X"FD",
X"F8",
X"F4",
X"F3",
X"F3",
X"F4",
X"F3",
X"F2",
X"F5",
X"F8",
X"F9",
X"FB",
X"FE",
X"FF",
X"FE",
X"FD",
X"FD",
X"FF",
X"00",
X"01",
X"02",
X"04",
X"06",
X"07",
X"04",
X"01",
X"00",
X"FD",
X"FC",
X"F8",
X"F4",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F5",
X"F9",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"04",
X"05",
X"05",
X"04",
X"01",
X"02",
X"02",
X"04",
X"06",
X"06",
X"06",
X"05",
X"05",
X"06",
X"06",
X"05",
X"03",
X"03",
X"03",
X"01",
X"00",
X"FD",
X"FC",
X"FB",
X"FA",
X"F8",
X"F8",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FD",
X"FE",
X"00",
X"02",
X"05",
X"07",
X"09",
X"09",
X"08",
X"07",
X"07",
X"07",
X"08",
X"09",
X"0A",
X"0A",
X"08",
X"07",
X"06",
X"05",
X"04",
X"04",
X"03",
X"01",
X"01",
X"00",
X"00",
X"FE",
X"FB",
X"F9",
X"F8",
X"F6",
X"F6",
X"F5",
X"F7",
X"FA",
X"FC",
X"FD",
X"00",
X"00",
X"00",
X"00",
X"04",
X"06",
X"08",
X"0B",
X"0B",
X"0B",
X"08",
X"06",
X"04",
X"02",
X"02",
X"02",
X"03",
X"04",
X"04",
X"05",
X"06",
X"07",
X"06",
X"03",
X"01",
X"00",
X"FF",
X"FB",
X"F9",
X"F7",
X"F6",
X"F4",
X"F3",
X"F3",
X"F2",
X"F3",
X"F5",
X"F6",
X"F6",
X"F7",
X"FA",
X"FD",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"04",
X"05",
X"06",
X"06",
X"05",
X"03",
X"01",
X"00",
X"FD",
X"FB",
X"F8",
X"F5",
X"F3",
X"F1",
X"EF",
X"EF",
X"EF",
X"EF",
X"F1",
X"F2",
X"F4",
X"F8",
X"FC",
X"00",
X"01",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"01",
X"01",
X"01",
X"03",
X"04",
X"04",
X"04",
X"05",
X"04",
X"03",
X"03",
X"03",
X"04",
X"06",
X"06",
X"05",
X"05",
X"05",
X"06",
X"08",
X"09",
X"09",
X"07",
X"05",
X"02",
X"00",
X"FF",
X"FD",
X"FC",
X"FA",
X"F9",
X"FA",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"FA",
X"FB",
X"FC",
X"FC",
X"FD",
X"FD",
X"FE",
X"FF",
X"00",
X"01",
X"04",
X"05",
X"06",
X"07",
X"08",
X"08",
X"09",
X"09",
X"0A",
X"0B",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0A",
X"09",
X"09",
X"08",
X"07",
X"05",
X"02",
X"00",
X"FF",
X"FD",
X"FB",
X"F9",
X"F7",
X"F6",
X"F5",
X"F4",
X"F4",
X"F5",
X"F4",
X"F4",
X"F6",
X"F8",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FE",
X"00",
X"04",
X"05",
X"06",
X"06",
X"05",
X"04",
X"02",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FE",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FC",
X"F7",
X"F5",
X"F2",
X"F1",
X"F0",
X"F0",
X"F0",
X"F1",
X"F2",
X"F1",
X"F1",
X"F2",
X"F4",
X"F6",
X"F8",
X"FA",
X"FC",
X"FD",
X"FE",
X"00",
X"03",
X"06",
X"08",
X"09",
X"0A",
X"0A",
X"09",
X"09",
X"07",
X"06",
X"05",
X"05",
X"06",
X"06",
X"06",
X"05",
X"04",
X"03",
X"03",
X"03",
X"04",
X"05",
X"05",
X"05",
X"05",
X"04",
X"02",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FD",
X"FC",
X"FB",
X"FA",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F8",
X"F9",
X"FA",
X"FC",
X"FC",
X"FE",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"01",
X"04",
X"06",
X"08",
X"08",
X"09",
X"09",
X"08",
X"06",
X"04",
X"03",
X"03",
X"03",
X"03",
X"04",
X"04",
X"05",
X"05",
X"04",
X"04",
X"04",
X"03",
X"02",
X"02",
X"03",
X"03",
X"03",
X"03",
X"04",
X"05",
X"05",
X"04",
X"04",
X"03",
X"03",
X"02",
X"01",
X"00",
X"FF",
X"FC",
X"FA",
X"F9",
X"F9",
X"F8",
X"F8",
X"F6",
X"F5",
X"F5",
X"F5",
X"F6",
X"F7",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FB",
X"FD",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"03",
X"04",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"06",
X"05",
X"05",
X"04",
X"02",
X"01",
X"00",
X"FF",
X"FD",
X"FC",
X"FA",
X"F8",
X"F7",
X"F5",
X"F4",
X"F2",
X"F2",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F5",
X"F7",
X"FA",
X"FC",
X"FF",
X"00",
X"01",
X"03",
X"04",
X"06",
X"06",
X"05",
X"05",
X"06",
X"06",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"03",
X"05",
X"06",
X"07",
X"08",
X"08",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"03",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FD",
X"FC",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"03",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"02",
X"02",
X"03",
X"03",
X"04",
X"04",
X"04",
X"06",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"05",
X"04",
X"03",
X"02",
X"01",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FA",
X"F9",
X"F8",
X"F7",
X"F6",
X"F5",
X"F4",
X"F3",
X"F2",
X"F1",
X"F1",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F3",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F7",
X"F8",
X"F9",
X"FA",
X"FB",
X"FB",
X"FC",
X"FE",
X"00",
X"00",
X"02",
X"03",
X"05",
X"07",
X"08",
X"09",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"08",
X"07",
X"06",
X"05",
X"05",
X"04",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"03",
X"03",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"04",
X"03",
X"03",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FB",
X"FB",
X"FA",
X"FA",
X"F9",
X"F9",
X"F8",
X"F8",
X"F7",
X"F7",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F9",
X"FA",
X"FA",
X"FB",
X"FD",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"02",
X"04",
X"05",
X"06",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"06",
X"06",
X"06",
X"06",
X"05",
X"05",
X"05",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"03",
X"02",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FB",
X"FA",
X"FA",
X"F8",
X"F7",
X"F6",
X"F5",
X"F3",
X"F2",
X"F2",
X"F1",
X"F1",
X"F1",
X"F0",
X"F0",
X"F0",
X"F1",
X"F2",
X"F2",
X"F3",
X"F4",
X"F5",
X"F6",
X"F7",
X"F8",
X"F9",
X"FA",
X"FB",
X"FC",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"01",
X"03",
X"03",
X"03",
X"05",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"04",
X"04",
X"04",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"02",
X"02",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"03",
X"03",
X"03",
X"04",
X"04",
X"04",
X"05",
X"05",
X"05",
X"05",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"02",
X"03",
X"03",
X"04",
X"04",
X"04",
X"05",
X"05",
X"05",
X"04",
X"04",
X"03",
X"03",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"02",
X"02",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"02",
X"03",
X"03",
X"04",
X"04",
X"05",
X"05",
X"05",
X"04",
X"04",
X"03",
X"03",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"03",
X"03",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FD",
X"FC",
X"FB",
X"FB",
X"FB",
X"FA",
X"FA",
X"FA",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FB",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"01",
X"01",
X"01",
X"02",
X"02",
X"02",
X"03",
X"04",
X"05",
X"05",
X"06",
X"06",
X"05",
X"04",
X"03",
X"02",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FC",
X"FC",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"FE",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"03",
X"04",
X"04",
X"05",
X"05",
X"04",
X"04",
X"03",
X"02",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"01",
X"01",
X"00",
X"00",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"02",
X"03",
X"03",
X"02",
X"01",
X"01",
X"00",
X"00",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FB",
X"FC",
X"FC",
X"FD",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FC",
X"FC",
X"FC",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"02",
X"03",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"02",
X"03",
X"04",
X"05",
X"06",
X"05",
X"04",
X"03",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FD",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FC",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"01",
X"02",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"03",
X"04",
X"04",
X"04",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FE",
X"FD",
X"FC",
X"FC",
X"FC",
X"FD",
X"FE",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FC",
X"FB",
X"FB",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FD",
X"FD",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"04",
X"04",
X"05",
X"05",
X"06",
X"05",
X"06",
X"06",
X"05",
X"04",
X"03",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FF",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FD",
X"FC",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"02",
X"02",
X"03",
X"04",
X"04",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"03",
X"01",
X"00",
X"FF",
X"FE",
X"FE",
X"FD",
X"FD",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"02",
X"03",
X"03",
X"04",
X"04",
X"03",
X"03",
X"03",
X"02",
X"02",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FD",
X"FC",
X"FB",
X"FA",
X"FA",
X"F9",
X"FA",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"02",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FE",
X"FE",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00"




  );
  begin

    if (RESET_N='0') then
      Q <= sin_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sin_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;