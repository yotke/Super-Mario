--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity coinTableTC is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(12 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end coinTableTC;

architecture arch of coinTableTC is

type table_type is array(0 to 8191) of std_logic_vector(7 downto 0);
signal sin_table : table_type;

begin

  SinTableTC_proc: process(RESET_N, CLK)
    constant sin_table : table_type := (
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"FD",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"04",
X"01",
X"FA",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"05",
X"04",
X"04",
X"03",
X"04",
X"03",
X"05",
X"FF",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"02",
X"05",
X"03",
X"04",
X"03",
X"04",
X"03",
X"05",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"01",
X"05",
X"03",
X"04",
X"03",
X"04",
X"03",
X"05",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"03",
X"04",
X"01",
X"FA",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"04",
X"03",
X"04",
X"03",
X"03",
X"04",
X"02",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"02",
X"05",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"01",
X"05",
X"03",
X"04",
X"03",
X"04",
X"03",
X"04",
X"FD",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"03",
X"04",
X"FE",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"03",
X"04",
X"02",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"FE",
X"05",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"04",
X"04",
X"03",
X"04",
X"03",
X"04",
X"03",
X"04",
X"FD",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"04",
X"03",
X"04",
X"03",
X"04",
X"03",
X"04",
X"FF",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FF",
X"05",
X"03",
X"04",
X"03",
X"03",
X"03",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FE",
X"04",
X"03",
X"04",
X"03",
X"03",
X"03",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FD",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"04",
X"01",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"02",
X"04",
X"03",
X"04",
X"03",
X"04",
X"02",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"02",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"02",
X"04",
X"01",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"01",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"FD",
X"FB",
X"FC",
X"FB",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"04",
X"FF",
X"FB",
X"FD",
X"FB",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"04",
X"00",
X"FA",
X"FD",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"FE",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"FE",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"04",
X"03",
X"03",
X"03",
X"03",
X"02",
X"04",
X"FF",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"02",
X"04",
X"03",
X"03",
X"03",
X"03",
X"02",
X"04",
X"00",
X"FB",
X"FD",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FE",
X"04",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"01",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"01",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"01",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FF",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FE",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FE",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"03",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"04",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"01",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"01",
X"FB",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"03",
X"02",
X"03",
X"02",
X"02",
X"03",
X"02",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"01",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"01",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FE",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"03",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"03",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FF",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"01",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"03",
X"01",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"01",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"03",
X"FF",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"FE",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"FF",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FF",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"01",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"01",
X"03",
X"02",
X"02",
X"02",
X"02",
X"01",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"01",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FF",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"00",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"00",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FF",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FD",
X"FD",
X"FD",
X"00",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"FE",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"05",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"01",
X"05",
X"03",
X"04",
X"03",
X"05",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"02",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FE",
X"05",
X"03",
X"04",
X"03",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"04",
X"04",
X"04",
X"04",
X"04",
X"02",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"02",
X"05",
X"03",
X"04",
X"03",
X"04",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"04",
X"04",
X"03",
X"04",
X"03",
X"04",
X"FE",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"02",
X"05",
X"03",
X"04",
X"03",
X"05",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"FE",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FF",
X"05",
X"03",
X"04",
X"03",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"04",
X"04",
X"04",
X"03",
X"04",
X"01",
X"FA",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"04",
X"03",
X"04",
X"04",
X"03",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"FE",
X"05",
X"04",
X"03",
X"03",
X"03",
X"04",
X"FD",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"04",
X"03",
X"04",
X"03",
X"04",
X"FF",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"01",
X"05",
X"03",
X"04",
X"03",
X"04",
X"FD",
X"FB",
X"FC",
X"FB",
X"FD",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"FF",
X"FA",
X"FC",
X"FB",
X"FD",
X"FB",
X"FF",
X"05",
X"03",
X"04",
X"03",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"01",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"FF",
X"05",
X"03",
X"04",
X"03",
X"03",
X"03",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FD",
X"04",
X"03",
X"03",
X"03",
X"04",
X"01",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"02",
X"04",
X"03",
X"03",
X"03",
X"03",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"04",
X"03",
X"04",
X"03",
X"04",
X"FE",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"02",
X"04",
X"03",
X"04",
X"02",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"02",
X"04",
X"02",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"05",
X"03",
X"04",
X"03",
X"04",
X"FF",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FE",
X"04",
X"03",
X"03",
X"03",
X"04",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FC",
X"FD",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"01",
X"04",
X"03",
X"03",
X"03",
X"03",
X"FD",
X"FB",
X"FC",
X"FC",
X"FC",
X"FD",
X"03",
X"03",
X"03",
X"03",
X"03",
X"04",
X"FE",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"02",
X"04",
X"02",
X"04",
X"02",
X"04",
X"00",
X"FB",
X"FC",
X"FB",
X"FD",
X"FB",
X"00",
X"04",
X"03",
X"03",
X"03",
X"04",
X"FE",
X"FB",
X"FD",
X"FB",
X"FD",
X"FB",
X"00",
X"04",
X"03",
X"03",
X"03",
X"04",
X"00",
X"FA",
X"FD",
X"FC",
X"FD",
X"FB",
X"FE",
X"04",
X"03",
X"03",
X"03",
X"04",
X"00",
X"FB",
X"FC",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FE",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"FD",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"01",
X"04",
X"03",
X"03",
X"03",
X"03",
X"FD",
X"FB",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"03",
X"03",
X"02",
X"04",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"01",
X"04",
X"02",
X"04",
X"02",
X"04",
X"00",
X"FB",
X"FC",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"02",
X"03",
X"02",
X"04",
X"01",
X"FB",
X"FC",
X"FC",
X"FD",
X"FC",
X"FF",
X"04",
X"02",
X"03",
X"02",
X"04",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"03",
X"03",
X"03",
X"03",
X"03",
X"01",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"02",
X"03",
X"03",
X"03",
X"03",
X"02",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"FE",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"02",
X"03",
X"02",
X"03",
X"02",
X"04",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"04",
X"00",
X"FB",
X"FC",
X"FC",
X"FD",
X"FB",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"04",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"03",
X"03",
X"03",
X"03",
X"03",
X"01",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FF",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"03",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FE",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"02",
X"03",
X"02",
X"03",
X"03",
X"02",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"FE",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"02",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FE",
X"04",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"02",
X"03",
X"03",
X"03",
X"03",
X"01",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"01",
X"03",
X"02",
X"03",
X"03",
X"03",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"01",
X"04",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"04",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"02",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FC",
X"FC",
X"FD",
X"FD",
X"FC",
X"FE",
X"03",
X"02",
X"02",
X"02",
X"02",
X"03",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"03",
X"02",
X"03",
X"FF",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"04",
X"02",
X"03",
X"02",
X"03",
X"01",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FE",
X"03",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"03",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"03",
X"02",
X"03",
X"01",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FF",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"03",
X"02",
X"02",
X"03",
X"01",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"01",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FE",
X"02",
X"03",
X"02",
X"02",
X"02",
X"03",
X"FF",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"01",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"03",
X"FF",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FE",
X"03",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FC",
X"FD",
X"FD",
X"FE",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FF",
X"FC",
X"FD",
X"FD",
X"FE",
X"FC",
X"FF",
X"03",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FF",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"03",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"01",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"02",
X"02",
X"02",
X"01",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"00",
X"03",
X"01",
X"02",
X"01",
X"03",
X"00",
X"FC",
X"FD",
X"FD",
X"FE",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"01",
X"03",
X"00",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"FF",
X"03",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FF",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FF",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"01",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FF",
X"FC",
X"FE",
X"FD",
X"FE",
X"FC",
X"00",
X"03",
X"02",
X"02",
X"01",
X"02",
X"00",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"FF",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FC",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"01",
X"02",
X"01",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FF",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"02",
X"02",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"01",
X"02",
X"01",
X"02",
X"FF",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"01",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"02",
X"02",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FD",
X"01",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FF",
X"02",
X"02",
X"02",
X"02",
X"01",
X"02",
X"FE",
X"FD",
X"FE",
X"FD",
X"FD",
X"FE",
X"01",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"FF",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"03",
X"01",
X"02",
X"01",
X"02",
X"01",
X"FE",
X"FD",
X"FE",
X"FE",
X"FD",
X"FE",
X"02",
X"02",
X"01",
X"02",
X"01",
X"02",
X"FF",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"01",
X"02",
X"01",
X"02",
X"02",
X"01",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"FF",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"01",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FF",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"01",
X"02",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"01",
X"FE",
X"FD",
X"FE",
X"FE",
X"FD",
X"FE",
X"02",
X"02",
X"01",
X"02",
X"01",
X"02",
X"FF",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"FF",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FF",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"FF",
X"02",
X"01",
X"01",
X"01",
X"01",
X"02",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"01",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"FF",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"02",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FF",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"FF",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"01",
X"01",
X"02",
X"FF",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"02",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"02",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FD",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FD",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"FF",
X"FE",
X"FF",
X"FE",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"01",
X"00",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FF",
X"FE",
X"FF",
X"FF",
X"FE",
X"FF",
X"01",
X"01",
X"00",
X"01",
X"00",
X"01",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"FF",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"01",
X"00",
X"00",
X"00",
X"00",
X"01",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00"







  );
  begin

    if (RESET_N='0') then
      Q <= sin_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sin_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;