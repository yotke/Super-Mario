library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
-- Alex Grinshpun April 2017

entity pipe_object is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) ;
		keepflag    : out std_logic
	);
end pipe_object;

architecture behav of pipe_object is 

constant object_X_size : integer := 100;
constant object_Y_size : integer := 184;
constant R_high		: integer := 7;
constant R_low		: integer := 5;
constant G_high		: integer := 4;
constant G_low		: integer := 2;
constant B_high		: integer := 1;
constant B_low		: integer := 0;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"31", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"35", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"79", x"79", x"79", x"7D", x"7D", x"7D", x"9E", x"9E", x"9E", x"9E", x"9E", x"9E", x"BE", x"BE", x"BE", x"BE", x"BF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BF", x"BE", x"BE", x"BE", x"BE", x"BE", x"9E", x"9E", x"9E", x"9E", x"9E", x"7E", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59"),
(x"55", x"55", x"59", x"59", x"55", x"55", x"55", x"55", x"55", x"55", x"35", x"31", x"31", x"31", x"30", x"30", x"30", x"30", x"30", x"30", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"55", x"55", x"59", x"59", x"59", x"59", x"79", x"79", x"79", x"79", x"7D", x"7E", x"9E", x"9E", x"9E", x"9E", x"BE", x"BE", x"BE", x"BE", x"BE", x"BF", x"BF", x"BF", x"DF", x"DF", x"BF", x"BF", x"BF", x"BE", x"BE", x"BE", x"BE", x"9E", x"9E", x"9E", x"9E", x"9E", x"7E", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59"),
(x"59", x"59", x"55", x"35", x"31", x"2C", x"2C", x"0C", x"0C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"38", x"38", x"38", x"58", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"55", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"38", x"38", x"58", x"58", x"59"),
(x"55", x"55", x"35", x"31", x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"38"),
(x"2C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"10", x"10", x"10", x"10", x"30"),
(x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"08", x"08", x"08", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"08", x"0C", x"0C"),
(x"08", x"08", x"08", x"08", x"08", x"00", x"55", x"51", x"31", x"2C", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"2C", x"2C", x"00", x"08", x"08", x"08", x"08", x"08"),
(x"00", x"00", x"00", x"00", x"00", x"55", x"55", x"55", x"31", x"2C", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"30", x"30", x"30", x"30", x"2C", x"2C", x"2C", x"2C", x"2C", x"2C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"08", x"08", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"55", x"55", x"55", x"31", x"2C", x"0C", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"2C", x"2C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"2C", x"2C", x"2C", x"2C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"55", x"55", x"55", x"31", x"2C", x"2C", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"2C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"2C", x"2C", x"2C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"55", x"55", x"55", x"31", x"2C", x"2C", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"2C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"2C", x"2C", x"2C", x"2C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"55", x"55", x"35", x"31", x"2C", x"08", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"2C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"55", x"55", x"35", x"31", x"2C", x"0C", x"08", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"35", x"35", x"55", x"55", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"55", x"55", x"55", x"31", x"2C", x"0C", x"08", x"08", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"2C", x"30", x"30", x"30", x"34", x"35", x"55", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"55", x"55", x"31", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"34", x"34", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"55", x"55", x"31", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"55", x"55", x"31", x"30", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"04", x"04", x"04", x"04", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"0C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"59", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"38", x"38", x"58", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"38", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"7D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"7D", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"79", x"7D", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"5D", x"5D", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"55", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"38", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"59", x"59", x"59", x"55", x"31", x"30", x"2C", x"0C", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"2C", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"34", x"34", x"34", x"34", x"34", x"34", x"54", x"54", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"59", x"58", x"58", x"58", x"58", x"38", x"38", x"34", x"34", x"34", x"34", x"34", x"38", x"38", x"58", x"59", x"59", x"00", x"00", x"00", x"00", x"00")
);
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000")
);


signal bCoord_X : integer := 0;
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--		
signal objectWestXboundary : integer;
signal objectSouthboundary : integer;
signal objectXboundariesTrue : boolean;
signal objectYboundariesTrue : boolean;
signal ObjectStartX_d : integer;
--signal keepflag : std_logic;
attribute syn_keep: boolean;
attribute syn_keep of keepflag: signal is true;
attribute preserve : boolean;
attribute preserve of keepflag: signal is true;
attribute noprune: boolean;  
attribute noprune of keepflag: signal is true;
begin

-- Calculate object boundaries
objectWestXboundary	<= object_X_size+ObjectStartX;
objectSouthboundary	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectWestXboundary) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectSouthboundary) else '0';

	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)

  		
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;
		ObjectStartX_d <= 0;

		elsif CLK'event and CLK='1' then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
			ObjectStartX_d <= ObjectStartX;
	end if;

  end process;

	keepflag <= '1' when 	ObjectStartX - ObjectStartX_d > 100 else '0';	
		
end behav;		
		