--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SinTableTC is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(7 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end SinTableTC;

architecture arch of SinTableTC is

type table_type is array(0 to 255) of std_logic_vector(7 downto 0);
signal sin_table : table_type;

begin

  SinTableTC_proc: process(RESET_N, CLK)
    constant sin_table : table_type := (
X"7D",
X"7B",
X"79",
X"77",
X"75",
X"73",
X"71",
X"6F",
X"6D",
X"6B",
X"6A",
X"68",
X"66",
X"64",
X"62",
X"61",
X"5F",
X"5D",
X"5C",
X"5A",
X"58",
X"57",
X"55",
X"53",
X"52",
X"50",
X"4F",
X"4D",
X"4B",
X"4A",
X"48",
X"47",
X"45",
X"44",
X"43",
X"41",
X"40",
X"3E",
X"3D",
X"3C",
X"3A",
X"39",
X"38",
X"36",
X"35",
X"34",
X"32",
X"31",
X"30",
X"2F",
X"2D",
X"2C",
X"2B",
X"2A",
X"29",
X"28",
X"27",
X"25",
X"24",
X"23",
X"22",
X"21",
X"20",
X"1F",
X"1E",
X"1D",
X"1C",
X"1B",
X"1A",
X"1A",
X"19",
X"18",
X"17",
X"16",
X"15",
X"14",
X"14",
X"13",
X"12",
X"11",
X"11",
X"10",
X"0F",
X"0F",
X"0E",
X"0D",
X"0D",
X"0C",
X"0B",
X"0B",
X"0A",
X"0A",
X"09",
X"08",
X"08",
X"07",
X"07",
X"06",
X"06",
X"06",
X"05",
X"05",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"02",
X"02",
X"03",
X"03",
X"03",
X"04",
X"04",
X"04",
X"05",
X"05",
X"06",
X"06",
X"06",
X"07",
X"07",
X"08",
X"08",
X"09",
X"0A",
X"0A",
X"0B",
X"0B",
X"0C",
X"0D",
X"0D",
X"0E",
X"0F",
X"0F",
X"10",
X"11",
X"11",
X"12",
X"13",
X"14",
X"14",
X"15",
X"16",
X"17",
X"18",
X"19",
X"1A",
X"1A",
X"1B",
X"1C",
X"1D",
X"1E",
X"1F",
X"20",
X"21",
X"22",
X"23",
X"24",
X"25",
X"27",
X"28",
X"29",
X"2A",
X"2B",
X"2C",
X"2D",
X"2F",
X"30",
X"31",
X"32",
X"34",
X"35",
X"36",
X"38",
X"39",
X"3A",
X"3C",
X"3D",
X"3E",
X"40",
X"41",
X"43",
X"44",
X"45",
X"47",
X"48",
X"4A",
X"4B",
X"4D",
X"4F",
X"50",
X"52",
X"53",
X"55",
X"57",
X"58",
X"5A",
X"5C",
X"5D",
X"5F",
X"61",
X"62",
X"64",
X"66",
X"68",
X"6A",
X"6B",
X"6D",
X"6F",
X"71",
X"73",
X"75",
X"77",
X"79",
X"7B",
X"7D",
X"7F"
  );
  begin

    if (RESET_N='0') then
      Q <= sin_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sin_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;