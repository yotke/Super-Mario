library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
-- Alex Grinshpun April 2017

entity smileyface_object is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer range 0 to 700;
		oCoord_Y	: in integer range 0 to 700;
		ObjectStartX	: in integer range 0 to 700;
		ObjectStartY 	: in integer range 0 to 700;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) ;
		keepflag    : out std_logic
	);
end smileyface_object;

architecture behav of smileyface_object is 

constant object_X_size : integer := 63;
constant object_Y_size : integer := 63;
constant R_high		: integer := 7;
constant R_low		: integer := 5;
constant G_high		: integer := 4;
constant G_low		: integer := 2;
constant B_high		: integer := 1;
constant B_low		: integer := 0;

type ram_array is array(0 to object_X_size - 1 , 0 to object_Y_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ED", x"E0", x"E4", x"E4", x"E4", x"E4", x"E4", x"ED", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E9", x"E9", x"E4", x"E4", x"E4", x"E4", x"E4", x"E4", x"E4", x"E4", x"E4", x"F6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ED", x"E4", x"E4", x"E4", x"E4", x"E4", x"E4", x"E4", x"E9", x"E9", x"E9", x"E4", x"E4", x"E4", x"ED", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E9", x"E0", x"E4", x"E4", x"E4", x"E0", x"E0", x"E4", x"F2", x"FB", x"FB", x"F6", x"F2", x"E4", x"E4", x"E4", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ED", x"E4", x"E9", x"E4", x"E0", x"E0", x"E0", x"E0", x"E9", x"FF", x"F2", x"ED", x"E9", x"F6", x"ED", x"E4", x"40", x"E9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ED", x"E9", x"E9", x"E4", x"E0", x"E0", x"E0", x"E0", x"E4", x"E9", x"FB", x"ED", x"F2", x"F2", x"ED", x"ED", x"E4", x"E4", x"E4", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E9", x"E9", x"E4", x"E4", x"E0", x"E0", x"E0", x"E0", x"E0", x"C4", x"F6", x"ED", x"FB", x"FB", x"F2", x"E9", x"C0", x"E4", x"C0", x"E9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E9", x"FF", x"E9", x"E4", x"E0", x"E0", x"E0", x"C0", x"C0", x"C0", x"C0", x"C9", x"ED", x"E9", x"E5", x"E4", x"E4", x"E4", x"E4", x"E9", x"E8", x"E9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F2", x"E9", x"E9", x"C4", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", x"E0", x"E4", x"E4", x"E4", x"C4", x"C0", x"C0", x"C0", x"C0", x"C4", x"C4", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"CD", x"C8", x"C4", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", x"E4", x"E0", x"C0", x"A0", x"80", x"80", x"80", x"80", x"80", x"80", x"A0", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"C9", x"C4", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"E4", x"C0", x"A0", x"60", x"60", x"64", x"40", x"20", x"40", x"60", x"60", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"C4", x"C4", x"C4", x"C0", x"C0", x"C0", x"A0", x"A0", x"C4", x"C4", x"80", x"60", x"40", x"20", x"88", x"A9", x"68", x"88", x"88", x"60", x"60", x"80", x"60", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A4", x"C0", x"A4", x"A4", x"A0", x"A0", x"A0", x"A0", x"A4", x"A4", x"64", x"64", x"88", x"AD", x"AD", x"D1", x"F6", x"F6", x"F6", x"D6", x"CD", x"D1", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A4", x"A8", x"A4", x"A0", x"A0", x"A0", x"80", x"80", x"84", x"84", x"88", x"AD", x"D6", x"DB", x"FB", x"F6", x"FA", x"F6", x"92", x"DB", x"F6", x"FB", x"64", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A4", x"A4", x"80", x"80", x"80", x"60", x"40", x"44", x"88", x"AD", x"D1", x"F6", x"DB", x"4E", x"72", x"FA", x"FA", x"F6", x"49", x"B7", x"D6", x"64", x"64", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"84", x"40", x"80", x"60", x"40", x"40", x"40", x"44", x"AD", x"F6", x"F6", x"FA", x"96", x"25", x"2A", x"DB", x"FA", x"F6", x"B2", x"DB", x"DA", x"D6", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"A9", x"AD", x"AD", x"89", x"44", x"40", x"44", x"89", x"F6", x"F6", x"FA", x"B6", x"2E", x"4E", x"DB", x"F6", x"F6", x"FA", x"FF", x"FF", x"FF", x"FE", x"FF", x"FA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F5", x"F6", x"F5", x"D1", x"CD", x"AD", x"44", x"40", x"64", x"D1", x"F6", x"FA", x"FA", x"BB", x"BB", x"D6", x"D1", x"FA", x"FA", x"FF", x"FF", x"FF", x"FA", x"FA", x"FA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"D1", x"D1", x"F1", x"F1", x"D1", x"AD", x"64", x"44", x"68", x"D6", x"F6", x"AD", x"B1", x"D6", x"D6", x"AD", x"AD", x"F6", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"D1", x"AD", x"F1", x"F6", x"F1", x"D1", x"88", x"64", x"AD", x"F6", x"F6", x"68", x"24", x"44", x"48", x"44", x"89", x"D1", x"F6", x"FA", x"FA", x"F6", x"F5", x"B6", x"FA", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AD", x"F1", x"D1", x"F6", x"F6", x"F5", x"AD", x"88", x"D1", x"F6", x"FA", x"B1", x"44", x"24", x"24", x"24", x"24", x"68", x"AD", x"B1", x"AD", x"AD", x"AD", x"C8", x"FF", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AD", x"88", x"D1", x"F5", x"F1", x"D1", x"AD", x"D1", x"F6", x"F6", x"FA", x"F6", x"8D", x"24", x"24", x"24", x"00", x"24", x"24", x"68", x"D1", x"F1", x"6D", x"D6", x"FB", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A8", x"84", x"CD", x"AD", x"68", x"64", x"AD", x"D1", x"F6", x"F6", x"FA", x"F6", x"B1", x"B1", x"8D", x"44", x"68", x"8D", x"D1", x"F1", x"8D", x"49", x"92", x"FB", x"B6", x"B6", x"DB", x"DB", x"FF", x"FF", x"B2", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"20", x"20", x"64", x"AD", x"D1", x"D2", x"F6", x"F6", x"F6", x"F6", x"D6", x"D1", x"D1", x"F5", x"F1", x"CD", x"8D", x"6D", x"8E", x"B6", x"DB", x"92", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"20", x"00", x"20", x"64", x"89", x"AD", x"D1", x"D1", x"F6", x"F6", x"F6", x"F5", x"F5", x"D1", x"6E", x"FC", x"92", x"92", x"8E", x"92", x"92", x"6D", x"B6", x"DB", x"DB", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"ED", x"84", x"60", x"60", x"44", x"69", x"89", x"AD", x"D1", x"D5", x"D1", x"CD", x"85", x"2A", x"4F", x"ED", x"A4", x"8D", x"8E", x"92", x"92", x"92", x"B6", x"FF", x"DB", x"DB", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"C9", x"C4", x"C0", x"C0", x"C0", x"A0", x"45", x"06", x"29", x"49", x"64", x"84", x"A0", x"84", x"2A", x"72", x"D5", x"A0", x"85", x"92", x"92", x"B6", x"B6", x"B6", x"BB", x"B7", x"DB", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"CD", x"C4", x"E4", x"E0", x"E4", x"C0", x"C0", x"A0", x"26", x"0B", x"0B", x"46", x"65", x"46", x"2A", x"0B", x"2F", x"B5", x"A8", x"A0", x"89", x"B2", x"B6", x"B6", x"B6", x"B6", x"B7", x"B7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ED", x"DF", x"E4", x"E4", x"E4", x"E4", x"E4", x"E4", x"C0", x"C4", x"65", x"0A", x"4E", x"96", x"72", x"2B", x"2B", x"2B", x"0B", x"2E", x"85", x"A0", x"A0", x"84", x"B2", x"B6", x"B7", x"B6", x"B7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ED", x"E4", x"E9", x"E4", x"E0", x"E4", x"E4", x"E0", x"C0", x"C0", x"C0", x"84", x"26", x"95", x"FD", x"D9", x"4E", x"2B", x"2F", x"2F", x"0B", x"46", x"A0", x"A0", x"80", x"FF", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E9", x"E9", x"E4", x"E0", x"E4", x"E4", x"E0", x"C0", x"C0", x"C0", x"C0", x"65", x"0A", x"6D", x"D8", x"B5", x"4E", x"2F", x"2F", x"2F", x"2F", x"2A", x"85", x"A4", x"A0", x"A9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"E0", x"E4", x"E4", x"E4", x"E4", x"C0", x"C0", x"A4", x"A0", x"A0", x"80", x"2A", x"0B", x"2A", x"4E", x"2E", x"2F", x"2F", x"2F", x"2F", x"0F", x"2F", x"2F", x"2F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"C9", x"E4", x"E0", x"E4", x"E4", x"C0", x"84", x"84", x"80", x"65", x"2A", x"0B", x"0B", x"2B", x"2B", x"2B", x"2F", x"2F", x"2F", x"0F", x"0B", x"2B", x"2F", x"2F", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C4", x"C4", x"E4", x"E0", x"E4", x"C4", x"C4", x"25", x"25", x"26", x"0A", x"0A", x"0B", x"0B", x"2B", x"2B", x"2B", x"2B", x"2B", x"2B", x"0B", x"2B", x"2B", x"2F", x"2B", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C4", x"C4", x"C4", x"E0", x"E4", x"C4", x"C0", x"05", x"05", x"06", x"0A", x"0A", x"0A", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"2B", x"2F", x"2F", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C4", x"C4", x"C4", x"E0", x"E4", x"C0", x"A0", x"05", x"05", x"06", x"06", x"0A", x"0A", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"2B", x"4F", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C4", x"C4", x"C0", x"E4", x"E9", x"C5", x"A4", x"25", x"05", x"05", x"06", x"06", x"0A", x"0A", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0A", x"2A", x"2A", x"4F", x"4E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"C9", x"CD", x"CE", x"F6", x"FB", x"FB", x"DB", x"DB", x"05", x"05", x"06", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"2A", x"2A", x"2A", x"2A", x"4E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"05", x"06", x"06", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"2A", x"2A", x"2A", x"2A", x"06", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"DB", x"DB", x"DB", x"DB", x"FF", x"FF", x"FB", x"DB", x"4E", x"06", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"2A", x"2A", x"26", x"0A", x"0A", x"2B", x"73", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B7", x"B6", x"B7", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"BB", x"2A", x"06", x"0A", x"0A", x"0A", x"0A", x"06", x"05", x"05", x"05", x"06", x"0A", x"0A", x"2B", x"4F", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B7", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"72", x"06", x"0A", x"0A", x"0A", x"0A", x"06", x"00", x"05", x"06", x"06", x"0A", x"0A", x"2B", x"4F", x"2F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"00", x"DB", x"DF", x"FF", x"FF", x"FF", x"DB", x"DB", x"FF", x"92", x"06", x"0A", x"0A", x"0A", x"0A", x"05", x"01", x"05", x"06", x"06", x"0A", x"0A", x"2A", x"4E", x"2E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"DB", x"DB", x"DB", x"FF", x"FF", x"DB", x"DB", x"FF", x"B7", x"4A", x"0A", x"0A", x"0A", x"0A", x"0A", x"25", x"05", x"05", x"06", x"06", x"0A", x"0A", x"2A", x"4E", x"4E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"B6", x"B7", x"DB", x"DB", x"FF", x"FF", x"FF", x"DB", x"4E", x"06", x"0A", x"0A", x"0A", x"0A", x"0A", x"25", x"05", x"05", x"06", x"06", x"0A", x"0A", x"2A", x"02", x"4E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"DB", x"B7", x"DB", x"DB", x"DB", x"DB", x"FF", x"B7", x"2A", x"0A", x"0A", x"0A", x"0A", x"0A", x"2A", x"25", x"05", x"05", x"06", x"06", x"0A", x"0A", x"2A", x"2A", x"4E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"2A", x"2A", x"0A", x"0A", x"0A", x"0B", x"0A", x"2A", x"25", x"05", x"05", x"06", x"06", x"0A", x"2A", x"2A", x"4F", x"2B", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"DB", x"DB", x"B7", x"B6", x"06", x"2A", x"2A", x"0A", x"0A", x"0B", x"0A", x"0A", x"2A", x"05", x"05", x"05", x"06", x"06", x"0A", x"0A", x"2A", x"65", x"88", x"A8", x"A8", x"C8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2A", x"2A", x"2A", x"2A", x"0A", x"0A", x"0B", x"0A", x"0A", x"2A", x"05", x"05", x"05", x"06", x"06", x"0A", x"0A", x"2A", x"68", x"A8", x"A8", x"C8", x"A8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2A", x"25", x"2A", x"0A", x"0A", x"0A", x"0B", x"0A", x"0A", x"25", x"05", x"05", x"05", x"06", x"06", x"0A", x"26", x"44", x"88", x"A8", x"A8", x"A8", x"A8", x"A8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"26", x"25", x"2A", x"0A", x"0A", x"0A", x"0B", x"0A", x"0A", x"25", x"20", x"05", x"05", x"05", x"05", x"25", x"44", x"64", x"89", x"A8", x"A8", x"A8", x"A8", x"84", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"25", x"2A", x"0A", x"0A", x"0B", x"0B", x"0A", x"0A", x"25", x"40", x"40", x"20", x"20", x"40", x"40", x"44", x"64", x"88", x"88", x"84", x"84", x"84", x"84", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"25", x"26", x"2A", x"2A", x"2A", x"2A", x"0A", x"0A", x"2A", x"68", x"64", x"44", x"44", x"40", x"40", x"40", x"44", x"64", x"64", x"64", x"64", x"64", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"44", x"44", x"44", x"44", x"64", x"64", x"44", x"44", x"24", x"25", x"F9", x"AC", x"8C", x"68", x"44", x"64", x"44", x"44", x"44", x"68", x"88", x"F9", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"64", x"64", x"84", x"88", x"A8", x"A8", x"88", x"84", x"64", x"44", x"44", x"44", x"00", x"D1", x"D1", x"AD", x"AC", x"AC", x"AC", x"B1", x"D1", x"D1", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"64", x"64", x"84", x"A8", x"A8", x"A8", x"AC", x"A8", x"84", x"64", x"84", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"64", x"64", x"84", x"A8", x"A8", x"A8", x"AD", x"A8", x"84", x"64", x"84", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"44", x"44", x"64", x"84", x"A8", x"A8", x"A8", x"84", x"64", x"44", x"64", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"68", x"68", x"68", x"64", x"84", x"84", x"64", x"64", x"64", x"68", x"68", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"8D", x"B1", x"AD", x"AD", x"AC", x"8C", x"8C", x"AD", x"B1", x"F5", x"D1", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F5", x"D1", x"D5", x"D5", x"D5", x"D5", x"F5", x"F9", x"F5", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

type object_form is array (0 to object_X_size - 1 , 0 to object_Y_size - 1) of std_logic;
constant object : object_form := (
("000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000011111111000000000000000000000000000"),
("000000000000000000000000001111111111110000000000000000000000000"),
("000000000000000000000000111111111111111000000000000000000000000"),
("000000000000000000000001111111111111111000000000000000000000000"),
("000000000000000000000011111111111111111100000000000000000000000"),
("000000000000000000000111111111111111111100000000000000000000000"),
("000000000000000000000111111111111111111110000000000000000000000"),
("000000000000000000001111111111111111111111000000000000000000000"),
("000000000000000000011111111111111111111111100000000000000000000"),
("000000000000000000011111111111111111111111100000000000000000000"),
("000000000000000000011111111111111111111111100000000000000000000"),
("000000000000000000111111111111111111111111100000000000000000000"),
("000000000000000000111111111111111111111110000000000000000000000"),
("000000000000000000111111111111111111111110000000000000000000000"),
("000000000000000000111111111111111111111110000000000000000000000"),
("000000000000000000111111111111111111111111000000000000000000000"),
("000000000000000000111111111111111111111111100000000000000000000"),
("000000000000000000111111111111111111111111100000000000000000000"),
("000000000000000000111111111111111111111111111111100000000000000"),
("000000000000000000111111111111111111111111111111110000000000000"),
("000000000000000000111111111111111111111111111111111000000000000"),
("000000000000000000011111111111111110111111111111111000000000000"),
("000000000000000000001111111111111111111111111111111100000000000"),
("000000000000000000000011111111111111111111111111111100000000000"),
("000000000000000000000011101111111111111111111111111100000000000"),
("000000000000000000000000111111111111111111111111111100000000000"),
("000000000000000000000001111111111111111111111111111100000000000"),
("000000000000000000000011111111111111111111111111111000000000000"),
("000000000000000000000111111111111111111111111111110000000000000"),
("000000000000000000001111111111111111111111111110000000000000000"),
("000000000000000000001111111111111111111111111100000000000000000"),
("000000000000000000011111111111111111111111110000000000000000000"),
("000000000000000000011111111111111111111111111000000000000000000"),
("000000000000000000011111111111111111111111111000000000000000000"),
("000000000000000000011111111111111111111111111000000000000000000"),
("000000000000000000011111111111111111111111110000000000000000000"),
("000000000000000000011111111111111111111111110000000000000000000"),
("000000000000000000111111111111111111111111110000000000000000000"),
("000000000000000000111111111111111111111111110000000000000000000"),
("000000000000000000111111111111111111111111110000000000000000000"),
("000000000000000000111111111111111111111111110000000000000000000"),
("000000000000000000111111111111111110111111110000000000000000000"),
("000000000000000000101111111111111111111111110000000000000000000"),
("000000000000000000111111111111111111111111110000000000000000000"),
("000000000000000000111111111111111111111111110000000000000000000"),
("000000000000000000111111111111111111111111110000000000000000000"),
("000000000000000000011111111111111111111111110000000000000000000"),
("000000000000000000001111111111111111111111111110000000000000000"),
("000000000000000000000000111111111111111111111110000000000000000"),
("000000000000000000000000111111111111111111111111000000000000000"),
("000000000000000000000000111111111111111111111111000000000000000"),
("000000000000000000000000111111111111111111111111000000000000000"),
("000000000000000000000000111111111111111111111110000000000000000"),
("000000000000000000000000111111111111111111111110000000000000000"),
("000000000000000000000000111111111111011111111100000000000000000"),
("000000000000000000000000111111111111000000000000000000000000000"),
("000000000000000000000000111111111111000000000000000000000000000"),
("000000000000000000000000111111111111000000000000000000000000000"),
("000000000000000000000000111111111110000000000000000000000000000"),
("000000000000000000000000111111111110000000000000000000000000000"),
("000000000000000000000000011111111100000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000")
);



signal bCoord_X : integer := 0;
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--		
signal objectWestXboundary : integer;
signal objectSouthboundary : integer;
signal objectXboundariesTrue : boolean;
signal objectYboundariesTrue : boolean;
signal ObjectStartX_d : integer;
--signal keepflag : std_logic;
attribute syn_keep: boolean;
attribute syn_keep of keepflag: signal is true;
attribute preserve : boolean;
attribute preserve of keepflag: signal is true;
attribute noprune: boolean;  
attribute noprune of keepflag: signal is true;
begin

-- Calculate object boundaries
objectWestXboundary	<= object_X_size+ObjectStartX;
objectSouthboundary	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectWestXboundary) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectSouthboundary) else '0';

	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)

  		
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;
		ObjectStartX_d <= 0;

		elsif CLK'event and CLK='1' then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
			ObjectStartX_d <= ObjectStartX;
	end if;

  end process;

	keepflag <= '1' when 	ObjectStartX - ObjectStartX_d > 100 else '0';	
		
end behav;		
		